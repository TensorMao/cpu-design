`ifndef __DIVIDE_SV
`define __DIVIDE_SV
`ifdef VERILATOR

`else

`endif
module divide();
endmodule


`endif