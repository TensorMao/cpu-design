`ifndef __BR_SV
`define __BR_SV
`ifdef VERILATOR

`else

`endif
module br()
endmodule
`endif