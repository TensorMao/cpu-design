`ifndef __PARAM_SV
`define __PARAM_SV 
      `define ALUOP_WIDTH 5
`ifdef VERILATOR
  
`else
`endif

`endif