`ifndef __ALUBMUX_SV
`define __ALUBMUX_SV
`ifdef VERILATOR

`else


`endif
module alubmux(
    input [1:0]ALUB_M
    

);
endmodule

`endif